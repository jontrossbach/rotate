`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/07/2020 06:20:43 PM
// Design Name: 
// Module Name: circular_right_rotate
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module circular_right_rotate(
    input wire[31:0] a,
    input wire[31:0] b,
    output wire[31:0] o
    );
    
   
    assign o = b[4:0] == 'b00001 ? {a[1:0],a[31:2]}
              :b[4:0] == 'b00010 ? {a[2:0],a[31:3]}
              :b[4:0] == 'b00011 ? {a[3:0],a[31:4]}
              :b[4:0] == 'b00100 ? {a[4:0],a[31:5]}
              :b[4:0] == 'b00101 ? {a[5:0],a[31:6]}
              :b[4:0] == 'b00111 ? {a[6:0],a[31:7]}
              :b[4:0] == 'b01000 ? {a[7:0],a[31:8]}
              :b[4:0] == 'b01001 ? {a[8:0],a[31:9]}
              :b[4:0] == 'b01010 ? {a[9:0],a[31:10]}
              :b[4:0] == 'b01011 ? {a[10:0],a[31:11]}
              :b[4:0] == 'b01100 ? {a[11:0],a[31:12]}
              :b[4:0] == 'b01101 ? {a[12:0],a[31:13]}
              :b[4:0] == 'b01110 ? {a[13:0],a[31:14]}
              :b[4:0] == 'b01111 ? {a[14:0],a[31:15]}
              :b[4:0] == 'b10000 ? {a[15:0],a[31:16]}
              :b[4:0] == 'b10001 ? {a[16:0],a[31:17]}
              :b[4:0] == 'b10010 ? {a[17:0],a[31:18]}
              :b[4:0] == 'b10011 ? {a[18:0],a[31:19]}
              :b[4:0] == 'b10100 ? {a[19:0],a[31:20]}
              :b[4:0] == 'b10101 ? {a[20:0],a[31:21]}
              :b[4:0] == 'b10110 ? {a[21:0],a[31:22]}
              :b[4:0] == 'b10111 ? {a[22:0],a[31:23]}
              :b[4:0] == 'b11000 ? {a[23:0],a[31:24]}
              :b[4:0] == 'b11001 ? {a[24:0],a[31:25]}
              :b[4:0] == 'b11010 ? {a[25:0],a[31:26]}
              :b[4:0] == 'b11011 ? {a[26:0],a[31:27]}
              :b[4:0] == 'b11100 ? {a[27:0],a[31:28]}
              :b[4:0] == 'b11101 ? {a[28:0],a[31:29]}
              :b[4:0] == 'b11110 ? {a[29:0],a[31:30]}
              :b[4:0] == 'b11111 ? {a[30:0],a[31]}
              :a;
 endmodule
